`timescale 1ns/1ns
`include "q4.v"

module q4_tb();

reg a,b,c,d;
wire f;

q4 ins_q4(a,b,c,d,f);

initial
begin

$dumpfile("q4_tb.vcd");
$dumpvars(0,q4_tb);

a=0;b=0;c=0;d=0;
#10;
a=0;b=0;c=0;d=1;
#10;
a=0;b=0;c=1;d=0;
#10;
a=0;b=0;c=1;d=1;
#10;
a=0;b=1;c=0;d=0;
#10;
a=0;b=1;c=0;d=1;
#10;
a=0;b=1;c=1;d=0;
#10;
a=0;b=1;c=1;d=1;
#10;
a=1;b=0;c=0;d=0;
#10;
a=1;b=0;c=0;d=1;
#10;
a=1;b=0;c=1;d=0;
#10;
a=1;b=0;c=1;d=1;
#10;
a=1;b=1;c=0;d=0;
#10;
a=1;b=1;c=0;d=1;
#10;
a=1;b=1;c=1;d=0;
#10;
a=1;b=1;c=1;d=1;
#10;

end
endmodule